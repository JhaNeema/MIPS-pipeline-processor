bind EXEStage fpv_exestage fpv_model_exe(.*);
bind controller_verif fpv_controller fpv_model_cont(.*);
bind EXE_MEM_stages fpv_exememstage fpv_model_exemem(.*);
bind hazard_detection fpv_hazard fpv_model_hdu(.*);
//bind MIPS_Processor assertions_pipeline fpv_model(clk, rst, forward_EN);

