bind EXEStage fpv_exestage fpv_model_exe(.*);
bind controller_verif fpv_controller fpv_model_cont(.*);
bind MIPS_Processor fpv_stages fpv_model_mips(.*);
bind hazard_detection fpv_hazard fpv_model_hdu(.*);

