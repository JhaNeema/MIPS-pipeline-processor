bind controller_non_combo fpv_controller fpv_model_cont(.*);
bind hazard_detection fpv_hazard fpv_model_hdu(.*);
bind EXEStage fpv_exestage fpv_model_exe(.*);
bind MIPS_Processor fpv_stages fpv_model_mips(.*);