bind IFStage assertions check1(clk, rst, freeze, brTaken, brOffset, instruction, PC);

